-- Author : YeN7zM  2025/06/12
-- This project is for 2025 DSD_Fianl_Question3
-- Propose : Display the "KIRBY" provided by TA, you have to display it like a traffic light, ex. RED -> YELLOW -> GREEN
-- and them have to turn on and off in 3, 2 ,4 secs, respectively
-- Scoring: 20/40 (Only finised the static traffic light)
-- Final Score: 100 / 120 (99 (A+) in final grade, 1/35)
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Final_Q1 is port(
    --VGA_sync
    CLOCK_50: IN std_logic;--記得除頻25
    KEY: IN std_logic_vector(1 downto 1);
    VGA_HS,VGA_VS: OUT std_logic;
    --rgb
    VGA_R, VGA_G, VGA_B:  out std_logic_vector(3 downto 0)
);
end ;

architecture a of Final_Q1 is
    --VGA_sync\rgb
    signal RESET: std_logic;
    signal video_on: std_logic;
    signal row, col: integer;--row_counter\col_counter
    signal CLK_25Mhz: std_logic;

    signal RGB: std_logic_vector(11 downto 0);

    component VGA_sync is
        port
        (	
            CLOCK,RESET: IN std_logic;
            HOR_SYN,VER_SYN,video_on: OUT std_logic;
            row_counter:out INTEGER RANGE 0 TO 524;
            col_counter:out INTEGER RANGE 0 TO 799
            ); 
	end component;

    component CLK_GEN is
        generic( divisor: integer := 50_000_000 ); 
        port 
        (	
            clock_in				: IN	STD_LOGIC;
            clock_out			: OUT	STD_LOGIC); 
    end component;

    type BITMAP is array(0 to 63) of std_logic_vector(0 to 127);--32col*16row (10*20放大)->320*320
    constant kirby: BITMAP := (--00=0 01=1 10=2 11=3
       "00000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            "00000000000000001111010101010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            "00000000000000110101010101010101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            "00000000000011010101010101010101011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            "00000000001101010101010101010101010111000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "00000000001101010101010101010101010111000000111111010101010101010101010111111100000000000000000000000000000000000000000000000000",
            "00000000110101010101010101010101010101111111010101010101010101010101010101010111110000000000000000000000000000000000000000000000",
            "00000000110101010101010101010101010111010101010101010101010101010101010101010101011111000000000000000000000000000000000000000000",
            "00000000110101010101010101010101011101010101010101010101010101010101010101010101010101110000000000000000000000000000000000000000",
            "00000000110101010101010101010101110101010101010101010101010101010101010101010101010101011111000000000000000000000000000000000000",
            "00000000110101010101010101010101010101010101010101010101010101010101010101010101010101010101110000000000000000000000000000000000",
            "00000000110101010101010101010101010101010101010101010101010101010101010101010101010101010101011111111111111111110000000000000000",
            "00000000110101010101010101010101010101010101010101010101010101010101111111010101010101010101010111010101010101011100000000000000",
            "00000000110101010101010101010101010101010101111111010101010101010111010111110101010101010101010101110101010101010111000000000000",
            "00000000110101010101010101010101010101010101110101110101010101010111010101110101010101010101010101011101010101010101110000000000",
            "00000000110101010101010101010101010101010111010101111101010101010111010101110101010101010101010101011101010101010101011100000000",
            "00000000110101010101010101010101010101010111010101011101010101010111010101111101010101010101010101010101010101010101011100000000",
            "00000000111101010101010101010101010101010111010101011101010101010111010101111101010101010101010101010101010101010101011100000000",
            "00000000001101010101010101010101010101010111110101111101010101010111111111111101010101010101010101010101010101010101011100000000",
            "00000000001101010101110101010101010101010111111111111101010101010111111111111101010101010101010101010101010101010101011100000000",
            "00000000001111010111010101010101010101010111111111111101010101010111111111111101010101010101010101010101010101010101011100000000",
            "00000000000011010111010101010101010101010111111111111101010101010111111111111101010101010101010101010101010101010101011100000000",
            "00000000000011010111010101010101010101010101111111111101010101010111111111111101010101010101010101010101110101010101110000000000",
            "00000000000000110111010101010101010101010101111111111101010101010101111111110101010110010101010101010101110101010101110000000000",
            "00000000000000111101010101010101010101010101111111111101010101010101111111110101011001100110010101010101011101010111000000000000",
            "00000000000000001101010101010101011001100101011111110101010101010101011111010101100110011001100101010101011101011111000000000000",
            "00000000000000001101010101010101100110011001010111010101010101010101010101010101011001100110010101010101011101111100000000000000",
            "00000000000000001101010101010110011001100101010101010101111111111111010101010101010101011001010101010101011111110000000000000000",
            "00000000000000001101010101010101100110010101010101010111101010101011010101010101010101010101010101010101111100000000000000000000",
            "00000000000000001101010101010101010101010101010101010111101010101011010101010101010101010101010101010101111100000000000000000000",
            "00000000000000001101010101010101010101010101010101010101111010101011010101010101010101010101010101111111110000000000000000000000",
            "00000000000000001101010101010101010101010101010101010101011110101101010101010101010101010111111111101010101100000000000000000000",
            "00000000000000001101010101010101010101010101010101010101010111110101010101010101010111111110101010101010101011000000000000000000",
            "00000000000000000011010101010101010101010101010101010101010101010101010101010101011110101010101010101010101010110000000000000000",
            "00000000000000000011010101010101010101010101010101010101010101010101010101010111111010101010101010101010101010101100000000000000",
            "00000000000000000011010101010101010101010101010101010101010101010101010101011110101010101010101010101010101010101100000000000000",
            "00000000000000000000110101010101010101010101010101010101010101010101010101111010101010101010101010101010101010101100000000000000",
            "00000000000000000000110101010101010101010101010101010101010101010101010111101010101010101010101010101010101010101100000000000000",
            "00000000000000000000001101010101010101010101010101010101010101010101011110101010101010101010101010101010101010101100000000000000",
            "00000000000000000000001111010101010101010101010101010101010101010101011110101010101010101010101010101010101010101100000000000000",
            "00000000000000000000000011010101010101010101010101010101010101010101111010101010101010101010101010101010101010101100000000000000",
            "00000000000000000000000011110101010101010101010101010101010101010101111010101010101010101010101010101010101010110000000000000000",
            "00000000000000000000000011101101010101010101010101010101010101010111101010101010101010101010101010101010101010110000000000000000",
            "00000000000000000000000011101011010101010101010101010101010101010111101010101010101010101010101010101010101011000000000000000000",
            "00000000000000000000000011101010110101010101010101010101010101010111101010101010101010101010101010101010101100000000000000000000",
            "00000000000000000000000011101010101111010101010101010101010101011110101010101010101010101010101010101010110000000000000000000000",
            "00000000000000000000000011101010101010111101010101010101010101011110101010101010101010101010101010101010110000000000000000000000",
            "00000000000000000000000000111010101010101011110101010101010101010111101010101010101010101010101010101011000000000000000000000000",
            "00000000000000000000000000111010101010101010101111111111010101010111101010101010101010101010101010101100000000000000000000000000",
            "00000000000000000000000000111010101010101010101010101010111111111111101010101010101010101010101010110000000000000000000000000000",
            "00000000000000000000000000111010101010101010101010101010101010101011111010101010101010101010101011000000000000000000000000000000",
            "00000000000000000000000000111010101010101010101010101010101010101011001110101010101010101010111100000000000000000000000000000000",
            "00000000000000000000000000001110101010101010101010101010101010101011001111101010101010101111000000000000000000000000000000000000",
            "00000000000000000000000000001110101010101010101010101010101010101011000000111111111111110000000000000000000000000000000000000000",
            "00000000000000000000000000001110101010101010101010101010101010101011000000000000000000000000000000000000000000000000000000000000",
            "00000000000000000000000000000011101010101010101010101010101010101011000000000000000000000000000000000000000000000000000000000000",
            "00000000000000000000000000000011101010101010101010101010101010101100000000000000000000000000000000000000000000000000000000000000",
            "00000000000000000000000000000000111010101010101010101010101010101100000000000000000000000000000000000000000000000000000000000000",
            "00000000000000000000000000000000001110101010101010101010101010101100000000000000000000000000000000000000000000000000000000000000",
            "00000000000000000000000000000000000011101010101010101010101010101100000000000000000000000000000000000000000000000000000000000000",
            "00000000000000000000000000000000000000111010101010101010101010110000000000000000000000000000000000000000000000000000000000000000",
            "00000000000000000000000000000000000000001111101010101010101011000000000000000000000000000000000000000000000000000000000000000000",
            "00000000000000000000000000000000000000000000111110101010111100000000000000000000000000000000000000000000000000000000000000000000",
            "00000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000"
    );
	 
    constant WHITE: std_logic_vector(11 downto 0) := x"FFF";
    constant BLACK: std_logic_vector(11 downto 0) := x"000";
    constant MOMO_PINK: std_logic_vector(11 downto 0) := x"F69";
    constant PINK: std_logic_vector(11 downto 0) := x"F9B";

begin
    RESET<=KEY(1);
    CLK_U1: CLK_GEN generic map(divisor => 2) port map(CLOCK_50, CLK_25Mhz);
    --VGA_sync
    VGA_sync_U1: VGA_sync port map(CLOCK => CLK_25Mhz,RESET=>KEY(1),HOR_SYN=>VGA_HS,VER_SYN=>VGA_VS,video_on=>video_on,row_counter=>row,col_counter=>col);

    process(video_on, row, col)
       variable kirby_row: std_logic_vector(0 to 127);
        --
        variable idx     : integer ;
        variable pattern : std_logic_vector(0 to 1);
    begin
        if(video_on = '0') then
            RGB <= BLACK;
        elsif(row >= 100 and row < 228 and col >= 20 and col < 148) then
            kirby_row := kirby((row-100)/ 2);
				idx:= ((col - 20)/ 2) * 2;
				pattern:= kirby_row(idx)&kirby_row(idx+1);
            case pattern is
                when "00" => RGB <= x"0AE";
                when "01" => RGB <= x"F03";
                when "10" => RGB <= x"F0A";
                when "11" => RGB <= x"501";
            end case;
		  elsif (row >= 100 and row < 228 and col >= 150 and col < 278) then
		  kirby_row := kirby((row-100)/ 2);
				idx:= ((col - 150)/ 2) * 2;
				pattern:= kirby_row(idx)&kirby_row(idx+1);
            case pattern is
                when "00" => RGB <= x"0AE";
                when "01" => RGB <= x"FD0";
                when "10" => RGB <= x"F10";
                when "11" => RGB <= x"440";
            end case;
				elsif (row >= 100 and row < 228 and col >= 278 and col < 406) then
		  kirby_row := kirby((row-100)/ 2);
				idx:= ((col - 278)/ 2) * 2;
				pattern:= kirby_row(idx)&kirby_row(idx+1);
            case pattern is
                when "00" => RGB <= x"0AE";
                when "01" => RGB <= x"7F2";
                when "10" => RGB <= x"D70";
                when "11" => RGB <= x"240";
            end case;
        else
            RGB <= x"0AE";
        end if;
    end process;
    VGA_R <= RGB(11 downto 8);
    VGA_G <= RGB(7 downto 4);
    VGA_B <= RGB(3 downto 0);
end architecture;

Library ieee;
use IEEE.STD_Logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-- Module Generates Video Sync Signals for Video Montor Interface
-- RGB and Sync outputs tie directly to monitor conector pins
ENTITY VGA_sync IS   
	PORT(
		CLOCK,RESET: IN std_logic;
		HOR_SYN,VER_SYN,video_on: OUT std_logic;
        row_counter:out INTEGER RANGE 0 TO 524;		
        col_counter:out INTEGER RANGE 0 TO 799	);
END VGA_sync ;

ARCHITECTURE arch OF VGA_sync IS
SIGNAL h_count: INTEGER RANGE 0 TO 799;			
SIGNAL v_count: INTEGER RANGE 0 TO 524;		
BEGIN

--Generate Horizontal and Vertical Timing Signals for Video Signal
-- 
--  Horiz_sync  ------------------------------------__________--------
--  h_count     0                 639              660      755      799
--
	PROCESS(CLOCK,RESET)   
	BEGIN				  						
     IF RESET = '0' THEN  h_count <=0;
     ELSIF CLOCK'EVENT AND CLOCK='1' THEN 
          IF h_count = 799 then h_count<=0;          
		  ELSE h_count <= h_count + 1;
     	  END IF;
     END IF;
	END PROCESS;

--  Vert_sync   ----------------------------------_______------------
--  v_count         0             479            493   494         524
--
   PROCESS(CLOCK,RESET)    
	BEGIN				  						
     IF RESET = '0' THEN v_count <=0;
     ELSIF CLOCK'EVENT AND CLOCK='1' THEN 
         IF h_count = 799 then 
			IF v_count = 524 THEN v_count <=0;
			ELSE v_count <= v_count+1;     
			END IF;
         END IF;
    END IF;
	END PROCESS;

--Generate Horizontal Sync Signal using h_count	
  PROCESS (h_count)  
    BEGIN
		IF h_count >=660 and h_count<=755 THEN HOR_SYN <= '0';
		ELSE  HOR_SYN <= '1';
		END IF;  	
  END PROCESS;
  
--Generate Vertical Sync Signal using v_count
   PROCESS (v_count)  
 	BEGIN
		IF (v_count >= 493 AND v_count <=494) THEN VER_SYN <= '0';
		ELSE VER_SYN <= '1';
		END IF;  	
	END PROCESS; 

-- Generate Video on Screen Signals for Pixel Data
-- Video on = 1 indicates pixel are being displayed
  process (h_count, v_count)  
	begin
		 IF v_count >=480 and v_count<=524 THEN video_on<='0';  
         ELSE 
			IF h_count >=640 and h_count<=799 THEN video_on<='0';
			ELSE video_on<='1';
			END IF;
     	END IF;
end process;

row_counter<=v_count;
col_counter<=h_count;

END arch;

--
-- Generate the user-specified clock signal (setting by divisor)
-- 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity CLK_GEN is
	generic( divisor: integer := 50_000_000 );
	port 
	(	
		clock_in				: IN	STD_LOGIC;
		clock_out			: OUT	STD_LOGIC); 
end CLK_GEN;

architecture arch of CLK_GEN is
	signal count: integer range 0 to divisor := 0;
	signal CLK_out: STD_LOGIC;
begin
	
	process(clock_in)
	begin
		IF clock_in'event and clock_in='1' THEN
			IF count <  divisor/2-1 THEN
				count <= count + 1;
			ELSE
				count <= 0;
				CLK_out <= NOT CLK_out;
			END IF;
		END IF;
		clock_out <= CLK_out;
	end process;
	
end arch;