LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Lab03_01 IS
    PORT (  SW : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
            HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6));
END Lab03_01;

ARCHITECTURE Structure OF Lab03_01 IS
    SIGNAL Sel : STD_LOGIC;
    SIGNAL W, X, Y, Z : STD_LOGIC;
BEGIN 
    PROCESS(SW)
    BEGIN    
        CASE SW IS --
                WHEN "00" => HEX0 <= "1000010"; 
                WHEN "01" => HEX0 <= "0110000"; 
                WHEN "10" => HEX0 <= "0000001"; 
                WHEN "11" => HEX0 <= "1111111"; 
                
            END CASE;
        END PROCESS;
END Structure;