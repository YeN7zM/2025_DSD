LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Lab02 IS
	PORT (	SW : IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
	        HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6));
END Lab02;

ARCHITECTURE Structure OF Lab02 IS
	SIGNAL Sel : STD_LOGIC;
	SIGNAL W, X, Y, Z : STD_LOGIC;
BEGIN 
	PROCESS(SW)
	BEGIN	
		CASE SW IS --
				WHEN "0000" => HEX0 <= "0000001"; 
				WHEN "0001" => HEX0 <= "1001111"; 
				WHEN "0010" => HEX0 <= "0010010"; 
				WHEN "0011" => HEX0 <= "0000110"; 
				WHEN "0100" => HEX0 <= "1001100"; 
				WHEN "0101" => HEX0 <= "0100100"; 
				WHEN "0110" => HEX0 <= "0100000"; 
				WHEN "0111" => HEX0 <= "0001111"; 
				WHEN "1000" => HEX0 <= "0000000"; 
				WHEN "1001" => HEX0 <= "0000100"; 
				WHEN "1010" => HEX0 <= "0001000"; 
				WHEN "1011" => HEX0 <= "1100000"; 
				WHEN "1100" => HEX0 <= "0110001"; 
				WHEN "1101" => HEX0 <= "1000010"; 
				WHEN "1110" => HEX0 <= "0110000"; 
				WHEN "1111" => HEX0 <= "0111000"; 
			END CASE;
		END PROCESS;
END Structure;


