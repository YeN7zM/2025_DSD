-- This project is for practicing the DSD_Fianl
-- Propose : Display your Student ID